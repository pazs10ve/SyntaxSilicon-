module and_gate(output y, input x1, input x2);
    assign y = x1 & x2;
endmodule