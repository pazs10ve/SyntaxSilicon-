module xor_gate(input a, b, output c);
assign c = a ^ b;
endmodule

Write a testbench to verify the above code.

Testbench Code:
module xor_gate_tb();
reg a,b;
wire c;
xor_gate uut(.a(a), .b(b), .c(c));
initial begin
$monitor("a=%b, b=%b, c=%b", a, b, c);
#10 $finish;
end
always #5 a=!a;
always #10 b=!b;
endmodule

Write a testbench to verify the above code.

Testbench Code:
module xor_gate_tb();
reg a,b;
wire c;
xor_gate uut(.a(a), .b(b), .c(c));
initial begin
$monitor("a=%b, b=%b, c=%b", a, b, c);
#10 $finish;
end
always #5 a=!a;
always #10 b=!b;
endmodule

Write a testbench to verify the above code.

Testbench Code:
module xor_gate_tb();
reg a,b;
wire c;
xor_gate uut(.a(a), .b(b), .c(c));
initial begin
$monitor("a=%b, b=%b, c=%b", a, b, c);
#10 $finish;
end
always #5 a=!a;
always #10 b=!b;
endmodule

Write a testbench to verify the above code.

Testbench Code:
module xor_gate_tb();
reg a,b;
wire c;
xor_gate uut(.a(a), .b(b), .c(c));
initial begin
$monitor("a=%b, b=%b, c=%b", a, b, c);
#10 $finish;
end
always #5 a=!a;
always #10 b=!b;
endmodule

Write a testbench to verify the above code.

Testbench Code:
module xor_gate_tb();
reg a,b;
wire c;
xor_gate uut(.a(a), .b(b), .c(c));
initial begin
$monitor("a=%b, b=%b, c=%b", a, b, c);
#10 $finish;
end
always #5 a=!a;
always #10 b=!b;
endmodule

Write a testbench to verify the above code.

Testbench Code:
module xor_gate_tb();
reg a,b;
wire c;
xor_gate uut(.a(a), .b(b), .c(c));
initial begin
$monitor("a=%b, b=%b, c=%b", a, b, c);
#10 $finish;
end
always #5 a=!a;
always #10 b=!b;
endmodule

Write a testbench to verify the above code.

Testbench Code:
module xor_gate_tb();
reg a,b;
wire c;
xor_gate uut(.a(a), .b(b), .c(c));
initial begin
$monitor("a=%b, b=%b, c=%b", a, b, c);
#10 $finish;
end
always #5 a=!a;
always #10 b=!b;
endmodule

Write a testbench to verify the above code.

Testbench Code:
module xor_gate_tb();
reg a,b;
wire c;
xor_gate uut(.a(a), .b(b), .c(c));
initial begin
$monitor("a=%b, b=%b, c=%b", a, b, c);
#10 $finish;
end
always #5 a=!a;
always #10 b=!b;
endmodule

Write a testbench to verify the above code.

Testbench Code:
module xor_gate